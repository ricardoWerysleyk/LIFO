library ieee;
use ieee.std_logic_1164.all;

entity demux_1x1_16 is
   port (entry: in std_logic;
			sel: in  std_logic_vector(3 downto 0);
         saida0, saida1, saida2, saida3, saida4, saida5: out std_logic;
			saida6, saida7, saida8, saida9, saida10: out std_logic;
			saida11, saida12, saida13, saida14, saida15: out std_logic);
end demux_1x1_16;

architecture logica of demux_1x1_16 is
	begin
		process (sel, entry)
			begin
				case sel is
					when "0000" => 
					saida0 <= entry;
					saida1 <= '0';
					saida2 <= '0';
					saida3 <= '0';
					saida4 <= '0';
					saida5 <= '0';
					saida6 <= '0';
					saida7 <= '0';
					saida8 <= '0';
					saida9 <= '0';
					saida10 <= '0';
					saida11 <= '0';
					saida12 <= '0';
					saida13 <= '0';
					saida14 <= '0';
					saida15 <= '0';
					when "0001" =>
					saida0 <= '0';
					saida1 <= entry;
					saida2 <= '0';
					saida3 <= '0';
					saida4 <= '0';
					saida5 <= '0';
					saida6 <= '0';
					saida7 <= '0';
					saida8 <= '0';
					saida9 <= '0';
					saida10 <= '0';
					saida11 <= '0';
					saida12 <= '0';
					saida13 <= '0';
					saida14 <= '0';
					saida15 <= '0';
					when "0010" => 
					saida0 <= '0';
					saida1 <= '0';
					saida2 <= entry;
					saida3 <= '0';
					saida4 <= '0';
					saida5 <= '0';
					saida6 <= '0';
					saida7 <= '0';
					saida8 <= '0';
					saida9 <= '0';
					saida10 <= '0';
					saida11 <= '0';
					saida12 <= '0';
					saida13 <= '0';
					saida14 <= '0';
					saida15 <= '0';
					when "0011" => 
					saida0 <= '0';
					saida1 <= '0';
					saida2 <= '0';
					saida3 <= entry;
					saida4 <= '0';
					saida5 <= '0';
					saida6 <= '0';
					saida7 <= '0';
					saida8 <= '0';
					saida9 <= '0';
					saida10 <= '0';
					saida11 <= '0';
					saida12 <= '0';
					saida13 <= '0';
					saida14 <= '0';
					saida15 <= '0';
					when "0100" => 
					saida0 <= '0';
					saida1 <= '0';
					saida2 <= '0';
					saida3 <= '0';
					saida4 <= entry;
					saida5 <= '0';
					saida6 <= '0';
					saida7 <= '0';
					saida8 <= '0';
					saida9 <= '0';
					saida10 <= '0';
					saida11 <= '0';
					saida12 <= '0';
					saida13 <= '0';
					saida14 <= '0';
					saida15 <= '0';
					when "0101" => 
					saida0 <= '0';
					saida1 <= '0';
					saida2 <= '0';
					saida3 <= '0';
					saida4 <= '0';
					saida5 <= entry;
					saida6 <= '0';
					saida7 <= '0';
					saida8 <= '0';
					saida9 <= '0';
					saida10 <= '0';
					saida11 <= '0';
					saida12 <= '0';
					saida13 <= '0';
					saida14 <= '0';
					saida15 <= '0';
					when "0110" => 
					saida0 <= '0';
					saida1 <= '0';
					saida2 <= '0';
					saida3 <= '0';
					saida4 <= '0';
					saida5 <= '0';
					saida6 <= entry;
					saida7 <= '0';
					saida8 <= '0';
					saida9 <= '0';
					saida10 <= '0';
					saida11 <= '0';
					saida12 <= '0';
					saida13 <= '0';
					saida14 <= '0';
					saida15 <= '0';
					when "0111" => 
					saida0 <= '0';
					saida1 <= '0';
					saida2 <= '0';
					saida3 <= '0';
					saida4 <= '0';
					saida5 <= '0';
					saida6 <= '0';
					saida7 <= entry;
					saida8 <= '0';
					saida9 <= '0';
					saida10 <= '0';
					saida11 <= '0';
					saida12 <= '0';
					saida13 <= '0';
					saida14 <= '0';
					saida15 <= '0';
					when "1000" => 
					saida0 <= '0';
					saida1 <= '0';
					saida2 <= '0';
					saida3 <= '0';
					saida4 <= '0';
					saida5 <= '0';
					saida6 <= '0';
					saida7 <= '0';
					saida8 <= entry;
					saida9 <= '0';
					saida10 <= '0';
					saida11 <= '0';
					saida12 <= '0';
					saida13 <= '0';
					saida14 <= '0';
					saida15 <= '0';
					when "1001" => 
					saida0 <= '0';
					saida1 <= '0';
					saida2 <= '0';
					saida3 <= '0';
					saida4 <= '0';
					saida5 <= '0';
					saida6 <= '0';
					saida7 <= '0';
					saida8 <= '0';
					saida9 <= entry;
					saida10 <= '0';
					saida11 <= '0';
					saida12 <= '0';
					saida13 <= '0';
					saida14 <= '0';
					saida15 <= '0';
					when "1010" => 
					saida0 <= '0';
					saida1 <= '0';
					saida2 <= '0';
					saida3 <= '0';
					saida4 <= '0';
					saida5 <= '0';
					saida6 <= '0';
					saida7 <= '0';
					saida8 <= '0';
					saida9 <= '0';
					saida10 <= entry;
					saida11 <= '0';
					saida12 <= '0';
					saida13 <= '0';
					saida14 <= '0';
					saida15 <= '0';
					when "1011" => 
					saida0 <= '0';
					saida1 <= '0';
					saida2 <= '0';
					saida3 <= '0';
					saida4 <= '0';
					saida5 <= '0';
					saida6 <= '0';
					saida7 <= '0';
					saida8 <= '0';
					saida9 <= '0';
					saida10 <= '0';
					saida11 <= entry;
					saida12 <= '0';
					saida13 <= '0';
					saida14 <= '0';
					saida15 <= '0';
					when "1100" =>
					saida0 <= '0';
					saida1 <= '0';
					saida2 <= '0';
					saida3 <= '0';
					saida4 <= '0';
					saida5 <= '0';
					saida6 <= '0';
					saida7 <= '0';
					saida8 <= '0';
					saida9 <= '0';
					saida10 <= '0';
					saida11 <= '0';
					saida12 <= entry;
					saida13 <= '0';
					saida14 <= '0';
					saida15 <= '0';
					when "1101" => 
					saida0 <= '0';
					saida1 <= '0';
					saida2 <= '0';
					saida3 <= '0';
					saida4 <= '0';
					saida5 <= '0';
					saida6 <= '0';
					saida7 <= '0';
					saida8 <= '0';
					saida9 <= '0';
					saida10 <= '0';
					saida11 <= '0';
					saida12 <= '0';
					saida13 <= entry;
					saida14 <= '0';
					saida15 <= '0';
					when "1110" => 
					saida0 <= '0';
					saida1 <= '0';
					saida2 <= '0';
					saida3 <= '0';
					saida4 <= '0';
					saida5 <= '0';
					saida6 <= '0';
					saida7 <= '0';
					saida8 <= '0';
					saida9 <= '0';
					saida10 <= '0';
					saida11 <= '0';
					saida12 <= '0';
					saida13 <= '0';
					saida14 <= entry;
					saida15 <= '0';
					when "1111" => 
					saida0 <= '0';
					saida1 <= '0';
					saida2 <= '0';
					saida3 <= '0';
					saida4 <= '0';
					saida5 <= '0';
					saida6 <= '0';
					saida7 <= '0';
					saida8 <= '0';
					saida9 <= '0';
					saida10 <= '0';
					saida11 <= '0';
					saida12 <= '0';
					saida13 <= '0';
					saida14 <= '0';
					saida15 <= entry;
				end case;
		end process;
end logica;